module frameBuffer(	input logic Clk, VGACLK, DrawEn,
					input logic DRAWX, DRAWY,
					input logic [1:0] playerDir,
					output R, G, B
					)

	logic [] frame;

endmodule